`define PARAMS_INIT_9 \
	.INIT_00(slice_init('h00)), \
	.INIT_01(slice_init('h01)), \
	.INIT_02(slice_init('h02)), \
	.INIT_03(slice_init('h03)), \
	.INIT_04(slice_init('h04)), \
	.INIT_05(slice_init('h05)), \
	.INIT_06(slice_init('h06)), \
	.INIT_07(slice_init('h07)), \
	.INIT_08(slice_init('h08)), \
	.INIT_09(slice_init('h09)), \
	.INIT_0A(slice_init('h0a)), \
	.INIT_0B(slice_init('h0b)), \
	.INIT_0C(slice_init('h0c)), \
	.INIT_0D(slice_init('h0d)), \
	.INIT_0E(slice_init('h0e)), \
	.INIT_0F(slice_init('h0f)), \
	.INIT_10(slice_init('h10)), \
	.INIT_11(slice_init('h11)), \
	.INIT_12(slice_init('h12)), \
	.INIT_13(slice_init('h13)), \
	.INIT_14(slice_init('h14)), \
	.INIT_15(slice_init('h15)), \
	.INIT_16(slice_init('h16)), \
	.INIT_17(slice_init('h17)), \
	.INIT_18(slice_init('h18)), \
	.INIT_19(slice_init('h19)), \
	.INIT_1A(slice_init('h1a)), \
	.INIT_1B(slice_init('h1b)), \
	.INIT_1C(slice_init('h1c)), \
	.INIT_1D(slice_init('h1d)), \
	.INIT_1E(slice_init('h1e)), \
	.INIT_1F(slice_init('h1f)),

`define PARAMS_INITP_9 \
	.INITP_00(slice_initp('h00)), \
	.INITP_01(slice_initp('h01)), \
	.INITP_02(slice_initp('h02)), \
	.INITP_03(slice_initp('h03)),

`define PARAMS_INIT_18 \
	.INIT_00(slice_init('h00)), \
	.INIT_01(slice_init('h01)), \
	.INIT_02(slice_init('h02)), \
	.INIT_03(slice_init('h03)), \
	.INIT_04(slice_init('h04)), \
	.INIT_05(slice_init('h05)), \
	.INIT_06(slice_init('h06)), \
	.INIT_07(slice_init('h07)), \
	.INIT_08(slice_init('h08)), \
	.INIT_09(slice_init('h09)), \
	.INIT_0A(slice_init('h0a)), \
	.INIT_0B(slice_init('h0b)), \
	.INIT_0C(slice_init('h0c)), \
	.INIT_0D(slice_init('h0d)), \
	.INIT_0E(slice_init('h0e)), \
	.INIT_0F(slice_init('h0f)), \
	.INIT_10(slice_init('h10)), \
	.INIT_11(slice_init('h11)), \
	.INIT_12(slice_init('h12)), \
	.INIT_13(slice_init('h13)), \
	.INIT_14(slice_init('h14)), \
	.INIT_15(slice_init('h15)), \
	.INIT_16(slice_init('h16)), \
	.INIT_17(slice_init('h17)), \
	.INIT_18(slice_init('h18)), \
	.INIT_19(slice_init('h19)), \
	.INIT_1A(slice_init('h1a)), \
	.INIT_1B(slice_init('h1b)), \
	.INIT_1C(slice_init('h1c)), \
	.INIT_1D(slice_init('h1d)), \
	.INIT_1E(slice_init('h1e)), \
	.INIT_1F(slice_init('h1f)), \
	.INIT_20(slice_init('h20)), \
	.INIT_21(slice_init('h21)), \
	.INIT_22(slice_init('h22)), \
	.INIT_23(slice_init('h23)), \
	.INIT_24(slice_init('h24)), \
	.INIT_25(slice_init('h25)), \
	.INIT_26(slice_init('h26)), \
	.INIT_27(slice_init('h27)), \
	.INIT_28(slice_init('h28)), \
	.INIT_29(slice_init('h29)), \
	.INIT_2A(slice_init('h2a)), \
	.INIT_2B(slice_init('h2b)), \
	.INIT_2C(slice_init('h2c)), \
	.INIT_2D(slice_init('h2d)), \
	.INIT_2E(slice_init('h2e)), \
	.INIT_2F(slice_init('h2f)), \
	.INIT_30(slice_init('h30)), \
	.INIT_31(slice_init('h31)), \
	.INIT_32(slice_init('h32)), \
	.INIT_33(slice_init('h33)), \
	.INIT_34(slice_init('h34)), \
	.INIT_35(slice_init('h35)), \
	.INIT_36(slice_init('h36)), \
	.INIT_37(slice_init('h37)), \
	.INIT_38(slice_init('h38)), \
	.INIT_39(slice_init('h39)), \
	.INIT_3A(slice_init('h3a)), \
	.INIT_3B(slice_init('h3b)), \
	.INIT_3C(slice_init('h3c)), \
	.INIT_3D(slice_init('h3d)), \
	.INIT_3E(slice_init('h3e)), \
	.INIT_3F(slice_init('h3f)),

`define PARAMS_INIT_18_U \
	.INIT_00(slice_init('h40)), \
	.INIT_01(slice_init('h41)), \
	.INIT_02(slice_init('h42)), \
	.INIT_03(slice_init('h43)), \
	.INIT_04(slice_init('h44)), \
	.INIT_05(slice_init('h45)), \
	.INIT_06(slice_init('h46)), \
	.INIT_07(slice_init('h47)), \
	.INIT_08(slice_init('h48)), \
	.INIT_09(slice_init('h49)), \
	.INIT_0A(slice_init('h4a)), \
	.INIT_0B(slice_init('h4b)), \
	.INIT_0C(slice_init('h4c)), \
	.INIT_0D(slice_init('h4d)), \
	.INIT_0E(slice_init('h4e)), \
	.INIT_0F(slice_init('h4f)), \
	.INIT_10(slice_init('h50)), \
	.INIT_11(slice_init('h51)), \
	.INIT_12(slice_init('h52)), \
	.INIT_13(slice_init('h53)), \
	.INIT_14(slice_init('h54)), \
	.INIT_15(slice_init('h55)), \
	.INIT_16(slice_init('h56)), \
	.INIT_17(slice_init('h57)), \
	.INIT_18(slice_init('h58)), \
	.INIT_19(slice_init('h59)), \
	.INIT_1A(slice_init('h5a)), \
	.INIT_1B(slice_init('h5b)), \
	.INIT_1C(slice_init('h5c)), \
	.INIT_1D(slice_init('h5d)), \
	.INIT_1E(slice_init('h5e)), \
	.INIT_1F(slice_init('h5f)), \
	.INIT_20(slice_init('h60)), \
	.INIT_21(slice_init('h61)), \
	.INIT_22(slice_init('h62)), \
	.INIT_23(slice_init('h63)), \
	.INIT_24(slice_init('h64)), \
	.INIT_25(slice_init('h65)), \
	.INIT_26(slice_init('h66)), \
	.INIT_27(slice_init('h67)), \
	.INIT_28(slice_init('h68)), \
	.INIT_29(slice_init('h69)), \
	.INIT_2A(slice_init('h6a)), \
	.INIT_2B(slice_init('h6b)), \
	.INIT_2C(slice_init('h6c)), \
	.INIT_2D(slice_init('h6d)), \
	.INIT_2E(slice_init('h6e)), \
	.INIT_2F(slice_init('h6f)), \
	.INIT_30(slice_init('h70)), \
	.INIT_31(slice_init('h71)), \
	.INIT_32(slice_init('h72)), \
	.INIT_33(slice_init('h73)), \
	.INIT_34(slice_init('h74)), \
	.INIT_35(slice_init('h75)), \
	.INIT_36(slice_init('h76)), \
	.INIT_37(slice_init('h77)), \
	.INIT_38(slice_init('h78)), \
	.INIT_39(slice_init('h79)), \
	.INIT_3A(slice_init('h7a)), \
	.INIT_3B(slice_init('h7b)), \
	.INIT_3C(slice_init('h7c)), \
	.INIT_3D(slice_init('h7d)), \
	.INIT_3E(slice_init('h7e)), \
	.INIT_3F(slice_init('h7f)),

`define PARAMS_INITP_18 \
	.INITP_00(slice_initp('h00)), \
	.INITP_01(slice_initp('h01)), \
	.INITP_02(slice_initp('h02)), \
	.INITP_03(slice_initp('h03)), \
	.INITP_04(slice_initp('h04)), \
	.INITP_05(slice_initp('h05)), \
	.INITP_06(slice_initp('h06)), \
	.INITP_07(slice_initp('h07)),

`define PARAMS_INIT_36 \
	.INIT_00(slice_init('h00)), \
	.INIT_01(slice_init('h01)), \
	.INIT_02(slice_init('h02)), \
	.INIT_03(slice_init('h03)), \
	.INIT_04(slice_init('h04)), \
	.INIT_05(slice_init('h05)), \
	.INIT_06(slice_init('h06)), \
	.INIT_07(slice_init('h07)), \
	.INIT_08(slice_init('h08)), \
	.INIT_09(slice_init('h09)), \
	.INIT_0A(slice_init('h0a)), \
	.INIT_0B(slice_init('h0b)), \
	.INIT_0C(slice_init('h0c)), \
	.INIT_0D(slice_init('h0d)), \
	.INIT_0E(slice_init('h0e)), \
	.INIT_0F(slice_init('h0f)), \
	.INIT_10(slice_init('h10)), \
	.INIT_11(slice_init('h11)), \
	.INIT_12(slice_init('h12)), \
	.INIT_13(slice_init('h13)), \
	.INIT_14(slice_init('h14)), \
	.INIT_15(slice_init('h15)), \
	.INIT_16(slice_init('h16)), \
	.INIT_17(slice_init('h17)), \
	.INIT_18(slice_init('h18)), \
	.INIT_19(slice_init('h19)), \
	.INIT_1A(slice_init('h1a)), \
	.INIT_1B(slice_init('h1b)), \
	.INIT_1C(slice_init('h1c)), \
	.INIT_1D(slice_init('h1d)), \
	.INIT_1E(slice_init('h1e)), \
	.INIT_1F(slice_init('h1f)), \
	.INIT_20(slice_init('h20)), \
	.INIT_21(slice_init('h21)), \
	.INIT_22(slice_init('h22)), \
	.INIT_23(slice_init('h23)), \
	.INIT_24(slice_init('h24)), \
	.INIT_25(slice_init('h25)), \
	.INIT_26(slice_init('h26)), \
	.INIT_27(slice_init('h27)), \
	.INIT_28(slice_init('h28)), \
	.INIT_29(slice_init('h29)), \
	.INIT_2A(slice_init('h2a)), \
	.INIT_2B(slice_init('h2b)), \
	.INIT_2C(slice_init('h2c)), \
	.INIT_2D(slice_init('h2d)), \
	.INIT_2E(slice_init('h2e)), \
	.INIT_2F(slice_init('h2f)), \
	.INIT_30(slice_init('h30)), \
	.INIT_31(slice_init('h31)), \
	.INIT_32(slice_init('h32)), \
	.INIT_33(slice_init('h33)), \
	.INIT_34(slice_init('h34)), \
	.INIT_35(slice_init('h35)), \
	.INIT_36(slice_init('h36)), \
	.INIT_37(slice_init('h37)), \
	.INIT_38(slice_init('h38)), \
	.INIT_39(slice_init('h39)), \
	.INIT_3A(slice_init('h3a)), \
	.INIT_3B(slice_init('h3b)), \
	.INIT_3C(slice_init('h3c)), \
	.INIT_3D(slice_init('h3d)), \
	.INIT_3E(slice_init('h3e)), \
	.INIT_3F(slice_init('h3f)), \
	.INIT_40(slice_init('h40)), \
	.INIT_41(slice_init('h41)), \
	.INIT_42(slice_init('h42)), \
	.INIT_43(slice_init('h43)), \
	.INIT_44(slice_init('h44)), \
	.INIT_45(slice_init('h45)), \
	.INIT_46(slice_init('h46)), \
	.INIT_47(slice_init('h47)), \
	.INIT_48(slice_init('h48)), \
	.INIT_49(slice_init('h49)), \
	.INIT_4A(slice_init('h4a)), \
	.INIT_4B(slice_init('h4b)), \
	.INIT_4C(slice_init('h4c)), \
	.INIT_4D(slice_init('h4d)), \
	.INIT_4E(slice_init('h4e)), \
	.INIT_4F(slice_init('h4f)), \
	.INIT_50(slice_init('h50)), \
	.INIT_51(slice_init('h51)), \
	.INIT_52(slice_init('h52)), \
	.INIT_53(slice_init('h53)), \
	.INIT_54(slice_init('h54)), \
	.INIT_55(slice_init('h55)), \
	.INIT_56(slice_init('h56)), \
	.INIT_57(slice_init('h57)), \
	.INIT_58(slice_init('h58)), \
	.INIT_59(slice_init('h59)), \
	.INIT_5A(slice_init('h5a)), \
	.INIT_5B(slice_init('h5b)), \
	.INIT_5C(slice_init('h5c)), \
	.INIT_5D(slice_init('h5d)), \
	.INIT_5E(slice_init('h5e)), \
	.INIT_5F(slice_init('h5f)), \
	.INIT_60(slice_init('h60)), \
	.INIT_61(slice_init('h61)), \
	.INIT_62(slice_init('h62)), \
	.INIT_63(slice_init('h63)), \
	.INIT_64(slice_init('h64)), \
	.INIT_65(slice_init('h65)), \
	.INIT_66(slice_init('h66)), \
	.INIT_67(slice_init('h67)), \
	.INIT_68(slice_init('h68)), \
	.INIT_69(slice_init('h69)), \
	.INIT_6A(slice_init('h6a)), \
	.INIT_6B(slice_init('h6b)), \
	.INIT_6C(slice_init('h6c)), \
	.INIT_6D(slice_init('h6d)), \
	.INIT_6E(slice_init('h6e)), \
	.INIT_6F(slice_init('h6f)), \
	.INIT_70(slice_init('h70)), \
	.INIT_71(slice_init('h71)), \
	.INIT_72(slice_init('h72)), \
	.INIT_73(slice_init('h73)), \
	.INIT_74(slice_init('h74)), \
	.INIT_75(slice_init('h75)), \
	.INIT_76(slice_init('h76)), \
	.INIT_77(slice_init('h77)), \
	.INIT_78(slice_init('h78)), \
	.INIT_79(slice_init('h79)), \
	.INIT_7A(slice_init('h7a)), \
	.INIT_7B(slice_init('h7b)), \
	.INIT_7C(slice_init('h7c)), \
	.INIT_7D(slice_init('h7d)), \
	.INIT_7E(slice_init('h7e)), \
	.INIT_7F(slice_init('h7f)),

`define PARAMS_INIT_36_U \
	.INIT_00(slice_init('h80)), \
	.INIT_01(slice_init('h81)), \
	.INIT_02(slice_init('h82)), \
	.INIT_03(slice_init('h83)), \
	.INIT_04(slice_init('h84)), \
	.INIT_05(slice_init('h85)), \
	.INIT_06(slice_init('h86)), \
	.INIT_07(slice_init('h87)), \
	.INIT_08(slice_init('h88)), \
	.INIT_09(slice_init('h89)), \
	.INIT_0A(slice_init('h8a)), \
	.INIT_0B(slice_init('h8b)), \
	.INIT_0C(slice_init('h8c)), \
	.INIT_0D(slice_init('h8d)), \
	.INIT_0E(slice_init('h8e)), \
	.INIT_0F(slice_init('h8f)), \
	.INIT_10(slice_init('h90)), \
	.INIT_11(slice_init('h91)), \
	.INIT_12(slice_init('h92)), \
	.INIT_13(slice_init('h93)), \
	.INIT_14(slice_init('h94)), \
	.INIT_15(slice_init('h95)), \
	.INIT_16(slice_init('h96)), \
	.INIT_17(slice_init('h97)), \
	.INIT_18(slice_init('h98)), \
	.INIT_19(slice_init('h99)), \
	.INIT_1A(slice_init('h9a)), \
	.INIT_1B(slice_init('h9b)), \
	.INIT_1C(slice_init('h9c)), \
	.INIT_1D(slice_init('h9d)), \
	.INIT_1E(slice_init('h9e)), \
	.INIT_1F(slice_init('h9f)), \
	.INIT_20(slice_init('ha0)), \
	.INIT_21(slice_init('ha1)), \
	.INIT_22(slice_init('ha2)), \
	.INIT_23(slice_init('ha3)), \
	.INIT_24(slice_init('ha4)), \
	.INIT_25(slice_init('ha5)), \
	.INIT_26(slice_init('ha6)), \
	.INIT_27(slice_init('ha7)), \
	.INIT_28(slice_init('ha8)), \
	.INIT_29(slice_init('ha9)), \
	.INIT_2A(slice_init('haa)), \
	.INIT_2B(slice_init('hab)), \
	.INIT_2C(slice_init('hac)), \
	.INIT_2D(slice_init('had)), \
	.INIT_2E(slice_init('hae)), \
	.INIT_2F(slice_init('haf)), \
	.INIT_30(slice_init('hb0)), \
	.INIT_31(slice_init('hb1)), \
	.INIT_32(slice_init('hb2)), \
	.INIT_33(slice_init('hb3)), \
	.INIT_34(slice_init('hb4)), \
	.INIT_35(slice_init('hb5)), \
	.INIT_36(slice_init('hb6)), \
	.INIT_37(slice_init('hb7)), \
	.INIT_38(slice_init('hb8)), \
	.INIT_39(slice_init('hb9)), \
	.INIT_3A(slice_init('hba)), \
	.INIT_3B(slice_init('hbb)), \
	.INIT_3C(slice_init('hbc)), \
	.INIT_3D(slice_init('hbd)), \
	.INIT_3E(slice_init('hbe)), \
	.INIT_3F(slice_init('hbf)), \
	.INIT_40(slice_init('hc0)), \
	.INIT_41(slice_init('hc1)), \
	.INIT_42(slice_init('hc2)), \
	.INIT_43(slice_init('hc3)), \
	.INIT_44(slice_init('hc4)), \
	.INIT_45(slice_init('hc5)), \
	.INIT_46(slice_init('hc6)), \
	.INIT_47(slice_init('hc7)), \
	.INIT_48(slice_init('hc8)), \
	.INIT_49(slice_init('hc9)), \
	.INIT_4A(slice_init('hca)), \
	.INIT_4B(slice_init('hcb)), \
	.INIT_4C(slice_init('hcc)), \
	.INIT_4D(slice_init('hcd)), \
	.INIT_4E(slice_init('hce)), \
	.INIT_4F(slice_init('hcf)), \
	.INIT_50(slice_init('hd0)), \
	.INIT_51(slice_init('hd1)), \
	.INIT_52(slice_init('hd2)), \
	.INIT_53(slice_init('hd3)), \
	.INIT_54(slice_init('hd4)), \
	.INIT_55(slice_init('hd5)), \
	.INIT_56(slice_init('hd6)), \
	.INIT_57(slice_init('hd7)), \
	.INIT_58(slice_init('hd8)), \
	.INIT_59(slice_init('hd9)), \
	.INIT_5A(slice_init('hda)), \
	.INIT_5B(slice_init('hdb)), \
	.INIT_5C(slice_init('hdc)), \
	.INIT_5D(slice_init('hdd)), \
	.INIT_5E(slice_init('hde)), \
	.INIT_5F(slice_init('hdf)), \
	.INIT_60(slice_init('he0)), \
	.INIT_61(slice_init('he1)), \
	.INIT_62(slice_init('he2)), \
	.INIT_63(slice_init('he3)), \
	.INIT_64(slice_init('he4)), \
	.INIT_65(slice_init('he5)), \
	.INIT_66(slice_init('he6)), \
	.INIT_67(slice_init('he7)), \
	.INIT_68(slice_init('he8)), \
	.INIT_69(slice_init('he9)), \
	.INIT_6A(slice_init('hea)), \
	.INIT_6B(slice_init('heb)), \
	.INIT_6C(slice_init('hec)), \
	.INIT_6D(slice_init('hed)), \
	.INIT_6E(slice_init('hee)), \
	.INIT_6F(slice_init('hef)), \
	.INIT_70(slice_init('hf0)), \
	.INIT_71(slice_init('hf1)), \
	.INIT_72(slice_init('hf2)), \
	.INIT_73(slice_init('hf3)), \
	.INIT_74(slice_init('hf4)), \
	.INIT_75(slice_init('hf5)), \
	.INIT_76(slice_init('hf6)), \
	.INIT_77(slice_init('hf7)), \
	.INIT_78(slice_init('hf8)), \
	.INIT_79(slice_init('hf9)), \
	.INIT_7A(slice_init('hfa)), \
	.INIT_7B(slice_init('hfb)), \
	.INIT_7C(slice_init('hfc)), \
	.INIT_7D(slice_init('hfd)), \
	.INIT_7E(slice_init('hfe)), \
	.INIT_7F(slice_init('hff)),

`define PARAMS_INITP_36 \
	.INITP_00(slice_initp('h00)), \
	.INITP_01(slice_initp('h01)), \
	.INITP_02(slice_initp('h02)), \
	.INITP_03(slice_initp('h03)), \
	.INITP_04(slice_initp('h04)), \
	.INITP_05(slice_initp('h05)), \
	.INITP_06(slice_initp('h06)), \
	.INITP_07(slice_initp('h07)), \
	.INITP_08(slice_initp('h08)), \
	.INITP_09(slice_initp('h09)), \
	.INITP_0A(slice_initp('h0a)), \
	.INITP_0B(slice_initp('h0b)), \
	.INITP_0C(slice_initp('h0c)), \
	.INITP_0D(slice_initp('h0d)), \
	.INITP_0E(slice_initp('h0e)), \
	.INITP_0F(slice_initp('h0f)),

`define MAKE_DO(do, dop, rdata) \
	wire [63:0] do; \
	wire [7:0] dop; \
	assign rdata = { \
		dop[7], \
		do[63:56], \
		dop[6], \
		do[55:48], \
		dop[5], \
		do[47:40], \
		dop[4], \
		do[39:32], \
		dop[3], \
		do[31:24], \
		dop[2], \
		do[23:16], \
		dop[1], \
		do[15:8], \
		dop[0], \
		do[7:0] \
	};

`define MAKE_DI(di, dip, wdata) \
	wire [63:0] di; \
	wire [7:0] dip; \
	assign { \
		dip[7], \
		di[63:56], \
		dip[6], \
		di[55:48], \
		dip[5], \
		di[47:40], \
		dip[4], \
		di[39:32], \
		dip[3], \
		di[31:24], \
		dip[2], \
		di[23:16], \
		dip[1], \
		di[15:8], \
		dip[0], \
		di[7:0] \
	} = wdata;

function [71:0] ival;
	input integer width;
	input [71:0] val;
	if (width == 72)
		ival = {
			val[71],
			val[62],
			val[53],
			val[44],
			val[35],
			val[26],
			val[17],
			val[8],
			val[70:63],
			val[61:54],
			val[52:45],
			val[43:36],
			val[34:27],
			val[25:18],
			val[16:9],
			val[7:0]
		};
	else if (width == 36)
		ival = {
			val[35],
			val[26],
			val[17],
			val[8],
			val[34:27],
			val[25:18],
			val[16:9],
			val[7:0]
		};
	else if (width == 18)
		ival = {
			val[17],
			val[8],
			val[16:9],
			val[7:0]
		};
	else
		ival = val;
endfunction

function [255:0] slice_init;
	input integer idx;
	integer i;
	for (i = 0; i < 32; i = i + 1)
		slice_init[i*8+:8] = INIT[(idx * 32 + i)*9+:8];
endfunction

function [255:0] slice_initp;
	input integer idx;
	integer i;
	for (i = 0; i < 256; i = i + 1)
		slice_initp[i] = INIT[(idx * 256 + i)*9+8];
endfunction
