module $__ICE40_SPRAM_ (...);

input PORT_A_CLK;
input PORT_A_CLK_EN;
input PORT_A_WR_EN;
input [3:0] PORT_A_WR_BE;
input [13:0] PORT_A_ADDR;
input [15:0] PORT_A_WR_DATA;
output [15:0] PORT_A_RD_DATA;

SB_SPRAM256KA _TECHMAP_REPLACE_ (
	.ADDRESS(PORT_A_ADDR),
	.DATAIN(PORT_A_WR_DATA),
	.MASKWREN(PORT_A_WR_BE),
	.WREN(PORT_A_WR_EN),
	.CHIPSELECT(PORT_A_CLK_EN),
	.CLOCK(PORT_A_CLK),
	.STANDBY(1'b0),
	.SLEEP(1'b0),
	.POWEROFF(1'b1),
	.DATAOUT(PORT_A_RD_DATA),
);

endmodule
